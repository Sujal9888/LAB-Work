LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY NAND_GATE_SUJAL IS
PORT(
	A: IN STD_LOGIC;
	B: IN STD_LOGIC;
	Y: OUT STD_LOGIC
	);
END NAND_GATE_SUJAL;
ARCHITECTURE Behavior of NAND_GATE_SUJAL IS

BEGIN
Y<= NOT (A AND B);
END Behavior;
