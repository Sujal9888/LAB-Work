LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY OR_GATE_SUJAL IS
PORT(
	A: IN STD_LOGIC;
	B: IN STD_LOGIC;
	Y: OUT STD_LOGIC
	);
END OR_GATE_SUJAL;
ARCHITECTURE Behavior of OR_GATE_SUJAL IS

BEGIN
Y<= A OR B;
END Behavior;
