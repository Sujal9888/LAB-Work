LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY XOR_GATE_SUJAL IS
PORT(
	A: IN STD_LOGIC;
	B: IN STD_LOGIC;
	Y: OUT STD_LOGIC
	);
END XOR_GATE_SUJAL;
ARCHITECTURE Behavior of XOR_GATE_SUJAL IS

BEGIN
Y<= A XOR B;
END Behavior;