LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY XNOR_GATE_SUJAL IS
PORT(
	A: IN STD_LOGIC;
	B: IN STD_LOGIC;
	Y: OUT STD_LOGIC
	);
END XNOR_GATE_SUJAL;
ARCHITECTURE Behavior of XNOR_GATE_SUJAL IS

BEGIN
Y<= NOT(A XOR B);
END Behavior;
