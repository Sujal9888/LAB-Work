LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY NOR_GATE_SUJAL IS
PORT(
	A: IN STD_LOGIC;
	B: IN STD_LOGIC;
	Y: OUT STD_LOGIC
	);
END NOR_GATE_SUJAL;
ARCHITECTURE Behavior of NOR_GATE_SUJAL IS

BEGIN
Y<= NOT (A OR B);
END Behavior;

