LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY AND_GATE_SUJAL IS
PORT(
	A: IN STD_LOGIC;
	B: IN STD_LOGIC;
	Y: OUT STD_LOGIC
	);
END AND_GATE_SUJAL;
ARCHITECTURE Behavior of AND_GATE_SUJAL IS

BEGIN
Y<= A AND B;
END Behavior;
